library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library work;
--use work.DadesRAM.ALL;

PACKAGE Programes is
--  TYPE memdata IS ARRAY (0 to m_size_real) of STD_LOGIC_VECTOR (n_data_real downto 0);
constant RAM_size	: integer := 2**5 - 1;
type MemoriaRAM is array (0 to RAM_size) of std_logic_vector (31 downto 0);


  CONSTANT programa2 : MemoriaRAM := ( 
	("00110100000001110000000001000000"), -- 0x00 ori $7, $0, 64        (0x34070040)
	("00110100000010000000000001001000"), -- 0x04 ori $8, $0, 72        (0x34080048)
	("00110100000010010000000001100000"), -- 0x08 ori $9, $0, 96        (0x34090060)
	("10001100111010100000000000000000"), -- 0x0C lw $10, 0($7)         (0x8CEA0000)
	("00000000000000000110000000100000"), -- 0x10 add $12, $0, $0       (0x00006020)
	("10001101000010110000000000000000"), -- 0x14 lw $11, 0($8)			  	(0x8D0B0000)
	("00000001011011000110000000100000"), -- 0x18 add $12, $11, $12     (0x016C6020)
	("00100001010010101111111111111111"), -- 0x1C addi $10, $10, -1     (0x214AFFFF) 
	("00100001000010000000000000000100"), -- 0x20 addi $8, $8, 4        (0x21080004)
	("00100001010010100000000000000000"), -- 0x1C addi $10, $10, 0  //actualitzem els flags abans del bgez
	("00000101101000011111111111111010"), -- 0x30 bgez $13, offset
	("10101101001011000000000000000000"), -- 0x34 sw $12, 0($9)         (0xAD2C0000)
	("00110100000010000000000000000010"), --  ori $8, $0, 2        (0x34080048)
	("00000001000001110100100000000110"), -- slrv $8, $7, $9 (rs/rt/rd)
	("00000000000000000000000000000000"), -- 0x30	              
	("00000000000000000000000000000000"), -- 0x34
	("00000000000000000000000000000000"), -- 0x38	
	("00000000000000000000000000000000"), -- 0x3C
	("00000000000000000000000000000101"), -- 0x40 5                     (0x00000005)
	("00000000000000000000000000000000"), -- 0x44 
	("00000000000000000000000101101101"), -- 0x48 365                   (0x0000016D)
	("00000000000000000000010111010100"), -- 0x4C 1492                  (0x000005D4)
	("00000000000000000000011111010001"), -- 0x50 2001                  (0x000007D1)
	("00000000000000000000001011000111"), -- 0x54 711                   (0x000002C7)
	("00000000000000000000011110011001"), -- 0x58 1945                  (0x00000799)
	("00000000000000000000000000000000"), -- 0x5C
	("00000000000000000000000000000000"), -- 0x60 0                     (0x00000000)
	("00000000000000000000000000000000"), -- 0x64
	("00000000000000000000000000000000"), -- 0x68
	("00000000000000000000000000000000"), -- 0x6C
	("00000000000000000000000000000000"), -- 
	("00000000000000000000000000000000") -- 0x70
  );

END Programes;